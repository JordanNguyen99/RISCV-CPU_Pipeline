��/ /  
 P h a s e  
 2  
 T e s t b e n c h  
 