��/ /  
 P h a s e  
 2  
 D a t a p a t h  
 