��m o d u l e   t e s t b e n c h ;  
  
         l o g i c   c l o c k ,   r e s e t ;  
         l o g i c   [ 3 1 : 0 ]   r e g i s t e r _ x 3 _ o u t ;  
  
         t o p   c p u _ t o p   (  
                 . c l o c k ( c l o c k ) ,  
                 . r e s e t ( r e s e t ) ,  
                 . r e g i s t e r _ x 3 _ o u t ( r e g i s t e r _ x 3 _ o u t )  
         ) ;  
  
         / /   C l o c k   g e n e r a t i o n  
         i n i t i a l   b e g i n  
                 c l o c k   =   0 ;  
                 f o r e v e r   # 5   c l o c k   =   ~ c l o c k ;   / /   C l o c k   p e r i o d   =   1 0   t i m e   u n i t s  
         e n d  
  
         / /   T e s t   s e q u e n c e  
         i n i t i a l   b e g i n  
                 r e s e t   =   1 ;  
                 # 1 0   r e s e t   =   0 ;  
  
                 # 1 0 0 ;  
                 $ d i s p l a y ( " R e g i s t e r   x 3   =   % 0 d " ,   r e g i s t e r _ x 3 _ o u t ) ;   / /   E x p e c t e d   o u t p u t :   1 5  
                 $ s t o p ;  
         e n d  
  
 e n d m o d u l e  
 