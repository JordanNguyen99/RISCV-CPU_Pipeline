��m o d u l e   d a t a p a t h   (  
         i n p u t     l o g i c   c l o c k ,                                   / /   S y s t e m   c l o c k  
         i n p u t     l o g i c   r e s e t ,                                   / /   A c t i v e - h i g h   r e s e t   s i g n a l  
         o u t p u t   l o g i c   [ 3 1 : 0 ]   r e g i s t e r _ x 3 _ o u t   / /   O u t p u t   r e g i s t e r   x 3   v a l u e   f o r   v e r i f i c a t i o n  
 ) ;  
  
         l o g i c   [ 3 1 : 0 ]   p r o g r a m _ c o u n t e r ,   n e x t _ p r o g r a m _ c o u n t e r ;  
         l o g i c   [ 3 1 : 0 ]   i n s t r u c t i o n ;  
         l o g i c   [ 3 1 : 0 ]   r e g i s t e r _ f i l e   [ 0 : 3 1 ] ;     / /   3 2   g e n e r a l - p u r p o s e   r e g i s t e r s  
  
         l o g i c   [ 3 1 : 0 ]   s o u r c e _ r e g i s t e r 1 _ d a t a ,   s o u r c e _ r e g i s t e r 2 _ d a t a ;  
         l o g i c   [ 3 1 : 0 ]   i m m e d i a t e _ v a l u e ;  
         l o g i c   [ 3 1 : 0 ]   a l u _ r e s u l t ;  
  
         l o g i c   [ 6 : 0 ]   o p c o d e ;  
         l o g i c   [ 4 : 0 ]   d e s t i n a t i o n _ r e g i s t e r ,   s o u r c e _ r e g i s t e r 1 ,   s o u r c e _ r e g i s t e r 2 ;  
         l o g i c   [ 2 : 0 ]   f u n c t 3 ;  
         l o g i c   [ 6 : 0 ]   f u n c t 7 ;  
  
         l o g i c   [ 3 1 : 0 ]   i n s t r u c t i o n _ m e m o r y   [ 0 : 1 5 ] ;   / /   H o l d s   p r o g r a m   i n s t r u c t i o n s  
  
         / /   L o a d   i n s t r u c t i o n s   f r o m   e x t e r n a l   f i l e   d u r i n g   s i m u l a t i o n  
         i n i t i a l   b e g i n  
                 $ r e a d m e m h ( " p r o g r a m . t x t " ,   i n s t r u c t i o n _ m e m o r y ) ;  
         e n d  
  
         / /   P r o g r a m   C o u n t e r   u p d a t e   l o g i c  
         a l w a y s _ f f   @ ( p o s e d g e   c l o c k   o r   p o s e d g e   r e s e t )   b e g i n  
                 i f   ( r e s e t )  
                         p r o g r a m _ c o u n t e r   < =   0 ;  
                 e l s e  
                         p r o g r a m _ c o u n t e r   < =   n e x t _ p r o g r a m _ c o u n t e r ;  
         e n d  
  
         a s s i g n   n e x t _ p r o g r a m _ c o u n t e r   =   p r o g r a m _ c o u n t e r   +   4 ;                               / /   W o r d - a l i g n e d  
         a s s i g n   i n s t r u c t i o n   =   i n s t r u c t i o n _ m e m o r y [ p r o g r a m _ c o u n t e r [ 5 : 2 ] ] ;     / /   F e t c h   i n s t r u c t i o n  
  
         / /   D e c o d e   i n s t r u c t i o n   f i e l d s  
         a s s i g n   o p c o d e   =   i n s t r u c t i o n [ 6 : 0 ] ;  
         a s s i g n   d e s t i n a t i o n _ r e g i s t e r   =   i n s t r u c t i o n [ 1 1 : 7 ] ;  
         a s s i g n   f u n c t 3   =   i n s t r u c t i o n [ 1 4 : 1 2 ] ;  
         a s s i g n   s o u r c e _ r e g i s t e r 1   =   i n s t r u c t i o n [ 1 9 : 1 5 ] ;  
         a s s i g n   s o u r c e _ r e g i s t e r 2   =   i n s t r u c t i o n [ 2 4 : 2 0 ] ;  
         a s s i g n   f u n c t 7   =   i n s t r u c t i o n [ 3 1 : 2 5 ] ;  
  
         / /   S i g n - e x t e n d   i m m e d i a t e   f o r   I - t y p e   i n s t r u c t i o n s  
         a s s i g n   i m m e d i a t e _ v a l u e   =   { { 2 0 { i n s t r u c t i o n [ 3 1 ] } } ,   i n s t r u c t i o n [ 3 1 : 2 0 ] } ;  
  
         / /   R e a d   r e g i s t e r   v a l u e s  
         a s s i g n   s o u r c e _ r e g i s t e r 1 _ d a t a   =   r e g i s t e r _ f i l e [ s o u r c e _ r e g i s t e r 1 ] ;  
         a s s i g n   s o u r c e _ r e g i s t e r 2 _ d a t a   =   r e g i s t e r _ f i l e [ s o u r c e _ r e g i s t e r 2 ] ;  
  
         / /   A L U   o p e r a t i o n :   s u p p o r t s   A D D I   a n d   A D D   i n s t r u c t i o n s  
         a s s i g n   a l u _ r e s u l t   =   ( o p c o d e   = =   7 ' b 0 0 1 0 0 1 1 )   ?   s o u r c e _ r e g i s t e r 1 _ d a t a   +   i m m e d i a t e _ v a l u e   :  
                                                 ( o p c o d e   = =   7 ' b 0 1 1 0 0 1 1 )   ?   s o u r c e _ r e g i s t e r 1 _ d a t a   +   s o u r c e _ r e g i s t e r 2 _ d a t a   :  
                                                 0 ;  
  
         / /   W r i t e   b a c k   r e s u l t   t o   d e s t i n a t i o n   r e g i s t e r  
         a l w a y s _ f f   @ ( p o s e d g e   c l o c k )   b e g i n  
                 i f   ( o p c o d e   = =   7 ' b 0 0 1 0 0 1 1   | |   o p c o d e   = =   7 ' b 0 1 1 0 0 1 1 )  
                         r e g i s t e r _ f i l e [ d e s t i n a t i o n _ r e g i s t e r ]   < =   a l u _ r e s u l t ;  
         e n d  
  
         / /   O u t p u t   r e g i s t e r   x 3   v a l u e  
         a s s i g n   r e g i s t e r _ x 3 _ o u t   =   r e g i s t e r _ f i l e [ 3 ] ;  
  
 e n d m o d u l e  
 