��/ /  
 P i p e l i n e  
 R e g i s t e r s  
 