��/ /  
 P h a s e  
 2  
 T o p  
 M o d u l e  
 