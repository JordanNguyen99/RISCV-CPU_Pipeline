��/ /  
 P h a s e  
 2  
 C o n t r o l  
 L o g i c  
 